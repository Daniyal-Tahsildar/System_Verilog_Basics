class common;
 static mailbox gen2drv_mbox = new();
 static semaphore smp = new(1);
endclass