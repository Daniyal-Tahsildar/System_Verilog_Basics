module queue;


endmodule