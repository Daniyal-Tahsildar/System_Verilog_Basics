interface intf (input logic clk);
    bit [5:0] ADDR, DATA, count;
endinterface