class common;
 static mailbox gen2drv_mbox = new();
endclass