class eth_common;
 static mailbox gen2bfm_mbox = new();

endclass